`timescale 1ns/1ps

module alu_test;

reg [31:0] instr;
reg signed [31:0] reg_A, reg_B;
wire signed [31:0] res;
wire [2:0] flags;

ALU testalu(instr, reg_A, reg_B, res, flags);

initial
begin

$display("instruction:op:func:   reg_A    :   reg_B    :   result   : flags");
$monitor("   %h:%h: %h :  %h  :  %h  :  %h  :  %h",
instr, testalu.opcode, testalu.func, testalu.regA, testalu.regB, testalu.result, testalu.flags);

#10 $display("add with no overflow");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;

#10 $display("add with possible overflow");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0000;
reg_A <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

#10 $display("addu");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0001;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0010_1000;

#10 $display("addu with possible overflow");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0001;
reg_A <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;
// flags = 0

#10 $display("Bitwise and");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0100;
reg_A <= 32'b0000_1100_0101_1001_0000_0110_1011_1100;
reg_B <= 32'b0000_0101_1001_1100_1000_1001_1001_0100;
// result: 32'b0000_0100_0001_1000_0000_0000_1001_0100(04180094 in hex)

#10 $display("Bitwise nor");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0111;
reg_A <= 32'b0011_1010_1111_0101_1100_0000_0001_1101;
reg_B <= 32'b0101_1010_0001_1100_1101_1000_0110_1001;
// result: 32'b1000_0101_0000_0010_0010_0111-1000_0010(85022782 in hex)

#10 $display("Bitwise or");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0101;
reg_A <= 32'b0000_1100_0101_1001_0000_0110_1011_1100;
reg_B <= 32'b0000_0101_1001_1100_1000_1001_1001_0100;
// result: 32'b0000_1101_1101_1101_1000_1111_1011_1100(0ddd8fbc in hex)

#10 $display("Shift left logical");
instr <= 32'b0000_0000_0000_0001_0000_0001_0000_0000;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
// result: 32'b0000_0000_0000_0000_0000_0010_0000_0000(00000200 in hex)

#10 $display("Shift left logical variable");
instr <= 32'b0000_0000_0000_0001_0000_0000_0000_0100;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
// result: 32'b0000_0000_0000_0000_0000_1000_0000_0000(00000800 in hex)

#10 $display("Set on less than with negative result");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_1010;
reg_A <= 32'b1000_0000_0000_0000_0000_0000_0001_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
// result: 32'b1, flag = 010(2 in hex)

#10 $display("Set on less than unsigned");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
reg_A <= 32'b1000_0000_0000_0000_0000_0000_0001_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
// flags = 000

#10 $display("Set on less than unsigned with negative result");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_1011;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
reg_B <= 32'b1000_0000_0000_0000_0000_0000_0010_0000;
// flags = 010(2 in hex)

#10 $display("Shift right arithmetic");
instr <= 32'b0000_0000_0000_0001_0000_0001_0000_0011;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
reg_B <= 32'b1000_0000_0000_0100_0000_0000_0000_0000;
// result: 32'b1111_1000_0000_0000_0100_0000_0000_0000(f8004000 in hex)

#10 $display("Shift right arithemetic variable");
instr <= 32'b0000_0000_0000_0001_0000_0000_0000_0111;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
reg_B <= 32'b1000_0000_1100_0100_0000_0000_0000_0000;
// result: 32'b1111_1111_1000_0000_1100_0100_0000_0000(ff80c400 in hex)

#10 $display("Shift right logical");
instr <= 32'b0000_0000_0000_0001_0000_0001_0000_0010;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
reg_B <= 32'b0000_1000_1100_0000_0000_0000_0000_0000;
// result: 32'b0000_0000_1000_1100_0000_0000_0000_0000(008c0000 in hex)

#10 $display("Shift right logical variable");
instr <= 32'b0000_0000_0000_0001_0000_0000_0000_0110;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
reg_B <= 32'b0000_1100_0011_0000_0000_0000_0000_0000;
// result: 32'b0000_0000_0000_1100_0011_0000_0000_0000(000c3000 in hex)

#10 $display("Subtract");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0010_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
// result: 32'b0000_0000_0000_0000_0000_0000_0001_1000(00000018 in hex)

#10 $display("Subtract with overflow");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0010;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg_B <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
// result: flag = 1

#10 $display("Subtract unsigned");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0011;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_0010;
reg_B <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;

#10 $display("Bitwise exclusive or");
instr <= 32'b0000_0000_0000_0001_0000_0000_0010_0110;
reg_A <= 32'b1001_0110_0011_1001_0010_0000_1111_0100;
reg_B <= 32'b0011_0100_1110_1101_0000_1010_0111_0000;
// result: 32'b1010_0010_1101_0100_0010_1010_1000_0100(a2d42a84 in hex)

#10 $display("Add immediate");
instr <= 32'b0010_0000_0000_0001_0000_0000_0011_0101;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0001_1100;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 32'b0000_0000_0000_0000_0000_0000_0101_0001(00000051 in hex)

#10 $display("Add immediate with overflow");
instr <= 32'b0010_0000_0000_0001_0000_0000_0011_0101;
reg_A <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 80000034 in hex  flag = 1

#10 $display("Add immediate unsigned");
instr <= 32'b0010_0100_0000_0001_0000_0000_0011_0101;
reg_A <= 32'b0111_1111_1111_1111_1111_1111_1111_1111;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 80000034 in hex  flag = 0

#10 $display("Branch on equal");
instr <= 32'b0001_0000_0000_0001_0000_0000_0000_1100;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1010;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1010;
// result: 00000030 flag = 4

#10 $display("Branch on not equal");
instr <= 32'b0001_0100_0000_0001_0000_0000_0000_1100;
reg_A <= 32'b0000_0000_0000_0000_0000_0000_0000_1010;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_1010;

#10 $display("Load word");
instr <= 32'b1000_1100_0000_0001_0000_0000_0000_0100;
reg_A <= 32'b0000_0000_0101_0000_0000_0000_0000_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 0x500004

#10 $display("Bitwise or immediate");
instr <= 32'b0011_0100_0000_0001_0011_1001_1100_0001;
reg_A <= 32'b0010_0011_1100_0000_1111_1110_0100_0101;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 32'b0010_0011_1100_0000_1111_1111_1100_0101(23c0ffc5 in hex)

#10 $display("Set on less than immediate");
instr <= 32'b0010_1000_0000_0001_1000_0000_0000_1010;
reg_A <= 32'b1111_1111_1111_1111_1000_0000_0000_1100;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

#10 $display("Set on less than immediate with negative result");
instr <= 32'b0010_1000_0000_0001_0000_0000_0000_1010;
reg_A <= 32'b1111_1111_1111_1111_1000_0000_0000_1001;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result:ffffffff      flags:010

#10 $display("Set on less than immediate unsigned");
instr <= 32'b0010_1100_0000_0001_1000_0000_0000_1010;
reg_A <= 32'b1111_1111_1111_1111_1000_0000_0000_1100;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

#10 $display("Set on less than immediate unsigned with negative result");
instr <= 32'b0010_1100_0000_0001_1000_0000_0000_1010;
reg_A <= 32'b1111_1111_1111_1111_1000_0000_0000_1001;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: ffffffff     flags: 010 

#10 $display("Store word");
instr <= 32'b1010_1100_0000_0001_0000_0000_0000_0100;
reg_A <= 32'b0000_0000_0101_0000_0000_0000_0000_0000;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;

#10 $display("Bitwise exclusive or immediate");
instr <= 32'b0011_1000_0000_0001_1110_0011_1010_0010;
reg_A <= 32'b0000_0110_1010_1000_0010_0101_1110_0001;
reg_B <= 32'b0000_0000_0000_0000_0000_0000_0000_0000;
// result: 32'b0000_0110_1010_1000_1100_0110_0100_0011(06a8c643 in hex)

#10 $finish;
end
endmodule